LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY ram IS
	PORT(
		clk : IN std_logic;
		we  : IN std_logic;
		address : IN  std_logic_vector(17 DOWNTO 0);
		datain  : IN  std_logic_vector(7 DOWNTO 0);
		dataout : OUT std_logic_vector(39 DOWNTO 0));
END ENTITY ram;

ARCHITECTURE syncrama OF ram IS

--64 kb Ram

	TYPE ram_type IS ARRAY(0 TO 262143) OF std_logic_vector(7 DOWNTO 0);
	SIGNAL ram : ram_type ;
	
	BEGIN
		PROCESS(clk) IS
			BEGIN
				IF rising_edge(clk) THEN  
					IF we = '1' THEN
						ram(to_integer(unsigned(address))) <= datain;
                                              
					END IF;
				END IF;
		END PROCESS;
--lower in lower and higher in higher
		dataout(7 downto 0) <= ram(to_integer(unsigned(address)));
                dataout(15 downto 8) <= ram(to_integer(unsigned(address))+1);
		dataout(23 downto 16) <= ram(to_integer(unsigned(address))+2);
		dataout(31 downto 24) <= ram(to_integer(unsigned(address))+3);
		dataout(39 downto 32) <= ram(to_integer(unsigned(address))+4);
END syncrama;
